module main

import utils

fn main() {
	println('Hello World!')

	println(utils.add(1, 2))
}
